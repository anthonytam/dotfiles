library verilog;
use verilog.vl_types.all;
entity Lab2 is
    port(
        \0\             : out    vl_logic;
        \1\             : out    vl_logic;
        \2\             : out    vl_logic;
        \3\             : out    vl_logic;
        \4\             : out    vl_logic;
        \5\             : out    vl_logic;
        \6\             : out    vl_logic;
        A               : in     vl_logic;
        C               : in     vl_logic;
        B               : in     vl_logic
    );
end Lab2;
